.param MOSFET_0_8_W_BIASCM_PMOS=2.0822112287558667 MOSFET_0_8_L_BIASCM_PMOS=0.6429299742183804 MOSFET_0_8_M_BIASCM_PMOS=27
.param MOSFET_8_2_W_gm1_PMOS=3.778524604683603 MOSFET_8_2_L_gm1_PMOS=0.2839144663858202 MOSFET_8_2_M_gm1_PMOS=77
.param MOSFET_10_1_W_gm2_PMOS=9.538962955988305 MOSFET_10_1_L_gm2_PMOS=0.8538902059252808 MOSFET_10_1_M_gm2_PMOS=22
.param MOSFET_11_1_W_gmf2_PMOS=8.36457886892506 MOSFET_11_1_L_gmf2_PMOS=0.15747933517957952 MOSFET_11_1_M_gmf2_PMOS=46
.param MOSFET_17_7_W_BIASCM_NMOS=1.6306712811825732 MOSFET_17_7_L_BIASCM_NMOS=0.7324691450349824 MOSFET_17_7_M_BIASCM_NMOS=47
.param MOSFET_21_2_W_LOAD2_NMOS=3.112627968762956 MOSFET_21_2_L_LOAD2_NMOS=0.7950677980821003 MOSFET_21_2_M_LOAD2_NMOS=92
.param MOSFET_23_1_W_gm3_NMOS=6.800388230019232 MOSFET_23_1_L_gm3_NMOS=0.7756911874818959 MOSFET_23_1_M_gm3_NMOS=2
.param CURRENT_0_BIAS=3.3724743993820217e-05
.param CAPACITOR_0=14.783740785188257e-12
.param CAPACITOR_1=92.81688379530945e-12
